** Profile: "SCHEMATIC1-Half"  [ C:\WORK\PROJECT\2_PLASMA_LF_GENERATOR\2_LF_GENERATOR_MAIN\4_REVIEW_DATA\Full_Bridge-PSpiceFiles\SCHEMATIC1\Half.sim ] 

** Creating circuit file "Half.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100us 0 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
