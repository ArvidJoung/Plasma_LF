** Profile: "SCHEMATIC1-LF_1stage"  [ E:\My_Work\20180114_Plasma_LF\2_LF_Generator_Main\4_Review_Data\lf_gen-pspicefiles\schematic1\lf_1stage.sim ] 

** Creating circuit file "LF_1stage.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100us 0 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
